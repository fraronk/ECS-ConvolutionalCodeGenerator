library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity CCG_tb is
    end entity CCG_tb;

    architecture bench of CCG_tb is

      constant T_CLK   : time := 8 ns;
      constant T_RESET : time := 15 ns;

        signal end_sim : std_logic := '1';
        signal clk_tb : std_logic := '0';
        signal rst_tb  : std_logic := '1';
        signal diff : std_logic;
        
        signal a_in_tb : std_logic;
        signal a_out_tb : std_logic;
        signal c_out_tb : std_logic;

        component CCG is
          port (
            clk : in std_logic;
            rst : in std_logic;
            a_in: in std_logic;
            a_out: out std_logic;
            c: out std_logic
          ) ;
        end component;

        signal t_integer : integer range 0 to 2047 := 0; -- t volte che si deve iterare il processo
        signal innp : std_logic_vector(10 downto 0) := "00000000000"; -- serie di 11 input che il dispositivo deve ricevere
        signal outp : std_logic_vector(10 downto 0) := "00000000000"; -- output calcolato passo passo
        signal count : std_logic_vector(11 downto 0) := "110000000000"; -- iteratore per tenere traccia al quale sottopasso siamo

        signal output_expected : std_logic_vector(10 downto 0); -- output aspettato al passo T
        type outp_t is array(natural range<>) of std_logic_vector(10 downto 0);
        -- la tabella sottostante contiene i risultati che si dovrebbero ottenere alla fine di ogni passo T, la tabella è stata generata dal codice java che simula il dispositivo
        constant outp_expected: outp_t := ("00000000000","10001100010","01000110001","11001010011","00100011000","10101111010","01100101001","11101001011","00010001100","10011101110","01010111101","11011011111","00110010100","10111110110","01110100101","11111000111","00001000110","10000100100","01001110111","11000010101","00101011110","10100111100","01101101111","11100001101","00011001010","10010101000","01011111011","11010011001","00111010010","10110110000","01111100011","11110000001","00000100011","10001000001","01000010010","11001110000","00100111011","10101011001","01100001010","11101101000","00010101111","10011001101","01010011110","11011111100","00110110111","10111010101","01110000110","11111100100","00001100101","10000000111","01001010100","11000110110","00101111101","10100011111","01101001100","11100101110","00011101001","10010001011","01011011000","11010111010","00111110001","10110010011","01111000000","11110100010","00000010001","10001110011","01000100000","11001000010","00100001001","10101101011","01100111000","11101011010","00010011101","10011111111","01010101100","11011001110","00110000101","10111100111","01110110100","11111010110","00001010111","10000110101","01001100110","11000000100","00101001111","10100101101","01101111110","11100011100","00011011011","10010111001","01011101010","11010001000","00111000011","10110100001","01111110010","11110010000","00000110010","10001010000","01000000011","11001100001","00100101010","10101001000","01100011011","11101111001","00010111110","10011011100","01010001111","11011101101","00110100110","10111000100","01110010111","11111110101","00001110100","10000010110","01001000101","11000100111","00101101100","10100001110","01101011101","11100111111","00011111000","10010011010","01011001001","11010101011","00111100000","10110000010","01111010001","11110110011","00000001000","10001101010","01000111001","11001011011","00100010000","10101110010","01100100001","11101000011","00010000100","10011100110","01010110101","11011010111","00110011100","10111111110","01110101101","11111001111","00001001110","10000101100","01001111111","11000011101","00101010110","10100110100","01101100111","11100000101","00011000010","10010100000","01011110011","11010010001","00111011010","10110111000","01111101011","11110001001","00000101011","10001001001","01000011010","11001111000","00100110011","10101010001","01100000010","11101100000","00010100111","10011000101","01010010110","11011110100","00110111111","10111011101","01110001110","11111101100","00001101101","10000001111","01001011100","11000111110","00101110101","10100010111","01101000100","11100100110","00011100001","10010000011","01011010000","11010110010","00111111001","10110011011","01111001000","11110101010","00000011001","10001111011","01000101000","11001001010","00100000001","10101100011","01100110000","11101010010","00010010101","10011110111","01010100100","11011000110","00110001101","10111101111","01110111100","11111011110","00001011111","10000111101","01001101110","11000001100","00101000111","10100100101","01101110110","11100010100","00011010011","10010110001","01011100010","11010000000","00111001011","10110101001","01111111010","11110011000","00000111010","10001011000","01000001011","11001101001","00100100010","10101000000","01100010011","11101110001","00010110110","10011010100","01010000111","11011100101","00110101110","10111001100","01110011111","11111111101","00001111100","10000011110","01001001101","11000101111","00101100100","10100000110","01101010101","11100110111","00011110000","10010010010","01011000001","11010100011","00111101000","10110001010","01111011001","11110111011","00000000100","10001100110","01000110101","11001010111","00100011100","10101111110","01100101101","11101001111","00010001000","10011101010","01010111001","11011011011","00110010000","10111110010","01110100001","11111000011","00001000010","10000100000","01001110011","11000010001","00101011010","10100111000","01101101011","11100001001","00011001110","10010101100","01011111111","11010011101","00111010110","10110110100","01111100111","11110000101","00000100111","10001000101","01000010110","11001110100","00100111111","10101011101","01100001110","11101101100","00010101011","10011001001","01010011010","11011111000","00110110011","10111010001","01110000010","11111100000","00001100001","10000000011","01001010000","11000110010","00101111001","10100011011","01101001000","11100101010","00011101101","10010001111","01011011100","11010111110","00111110101","10110010111","01111000100","11110100110","00000010101","10001110111","01000100100","11001000110","00100001101","10101101111","01100111100","11101011110","00010011001","10011111011","01010101000","11011001010","00110000001","10111100011","01110110000","11111010010","00001010011","10000110001","01001100010","11000000000","00101001011","10100101001","01101111010","11100011000","00011011111","10010111101","01011101110","11010001100","00111000111","10110100101","01111110110","11110010100","00000110110","10001010100","01000000111","11001100101","00100101110","10101001100","01100011111","11101111101","00010111010","10011011000","01010001011","11011101001","00110100010","10111000000","01110010011","11111110001","00001110000","10000010010","01001000001","11000100011","00101101000","10100001010","01101011001","11100111011","00011111100","10010011110","01011001101","11010101111","00111100100","10110000110","01111010101","11110110111","00000001100","10001101110","01000111101","11001011111","00100010100","10101110110","01100100101","11101000111","00010000000","10011100010","01010110001","11011010011","00110011000","10111111010","01110101001","11111001011","00001001010","10000101000","01001111011","11000011001","00101010010","10100110000","01101100011","11100000001","00011000110","10010100100","01011110111","11010010101","00111011110","10110111100","01111101111","11110001101","00000101111","10001001101","01000011110","11001111100","00100110111","10101010101","01100000110","11101100100","00010100011","10011000001","01010010010","11011110000","00110111011","10111011001","01110001010","11111101000","00001101001","10000001011","01001011000","11000111010","00101110001","10100010011","01101000000","11100100010","00011100101","10010000111","01011010100","11010110110","00111111101","10110011111","01111001100","11110101110","00000011101","10001111111","01000101100","11001001110","00100000101","10101100111","01100110100","11101010110","00010010001","10011110011","01010100000","11011000010","00110001001","10111101011","01110111000","11111011010","00001011011","10000111001","01001101010","11000001000","00101000011","10100100001","01101110010","11100010000","00011010111","10010110101","01011100110","11010000100","00111001111","10110101101","01111111110","11110011100","00000111110","10001011100","01000001111","11001101101","00100100110","10101000100","01100010111","11101110101","00010110010","10011010000","01010000011","11011100001","00110101010","10111001000","01110011011","11111111001","00001111000","10000011010","01001001001","11000101011","00101100000","10100000010","01101010001","11100110011","00011110100","10010010110","01011000101","11010100111","00111101100","10110001110","01111011101","11110111111","00000000010","10001100000","01000110011","11001010001","00100011010","10101111000","01100101011","11101001001","00010001110","10011101100","01010111111","11011011101","00110010110","10111110100","01110100111","11111000101","00001000100","10000100110","01001110101","11000010111","00101011100","10100111110","01101101101","11100001111","00011001000","10010101010","01011111001","11010011011","00111010000","10110110010","01111100001","11110000011","00000100001","10001000011","01000010000","11001110010","00100111001","10101011011","01100001000","11101101010","00010101101","10011001111","01010011100","11011111110","00110110101","10111010111","01110000100","11111100110","00001100111","10000000101","01001010110","11000110100","00101111111","10100011101","01101001110","11100101100","00011101011","10010001001","01011011010","11010111000","00111110011","10110010001","01111000010","11110100000","00000010011","10001110001","01000100010","11001000000","00100001011","10101101001","01100111010","11101011000","00010011111","10011111101","01010101110","11011001100","00110000111","10111100101","01110110110","11111010100","00001010101","10000110111","01001100100","11000000110","00101001101","10100101111","01101111100","11100011110","00011011001","10010111011","01011101000","11010001010","00111000001","10110100011","01111110000","11110010010","00000110000","10001010010","01000000001","11001100011","00100101000","10101001010","01100011001","11101111011","00010111100","10011011110","01010001101","11011101111","00110100100","10111000110","01110010101","11111110111","00001110110","10000010100","01001000111","11000100101","00101101110","10100001100","01101011111","11100111101","00011111010","10010011000","01011001011","11010101001","00111100010","10110000000","01111010011","11110110001","00000001010","10001101000","01000111011","11001011001","00100010010","10101110000","01100100011","11101000001","00010000110","10011100100","01010110111","11011010101","00110011110","10111111100","01110101111","11111001101","00001001100","10000101110","01001111101","11000011111","00101010100","10100110110","01101100101","11100000111","00011000000","10010100010","01011110001","11010010011","00111011000","10110111010","01111101001","11110001011","00000101001","10001001011","01000011000","11001111010","00100110001","10101010011","01100000000","11101100010","00010100101","10011000111","01010010100","11011110110","00110111101","10111011111","01110001100","11111101110","00001101111","10000001101","01001011110","11000111100","00101110111","10100010101","01101000110","11100100100","00011100011","10010000001","01011010010","11010110000","00111111011","10110011001","01111001010","11110101000","00000011011","10001111001","01000101010","11001001000","00100000011","10101100001","01100110010",
        "11101010000","00010010111","10011110101","01010100110","11011000100","00110001111","10111101101","01110111110","11111011100","00001011101","10000111111","01001101100","11000001110","00101000101","10100100111","01101110100","11100010110","00011010001","10010110011","01011100000","11010000010","00111001001","10110101011","01111111000","11110011010","00000111000","10001011010","01000001001","11001101011","00100100000","10101000010","01100010001","11101110011","00010110100","10011010110","01010000101","11011100111","00110101100","10111001110","01110011101","11111111111","00001111110","10000011100","01001001111","11000101101","00101100110","10100000100","01101010111","11100110101","00011110010","10010010000","01011000011","11010100001","00111101010","10110001000","01111011011","11110111001","00000000110","10001100100","01000110111","11001010101","00100011110","10101111100","01100101111","11101001101","00010001010","10011101000","01010111011","11011011001","00110010010","10111110000","01110100011","11111000001","00001000000","10000100010","01001110001","11000010011","00101011000","10100111010","01101101001","11100001011","00011001100","10010101110","01011111101","11010011111","00111010100","10110110110","01111100101","11110000111","00000100101","10001000111","01000010100","11001110110","00100111101","10101011111","01100001100","11101101110","00010101001","10011001011","01010011000","11011111010","00110110001","10111010011","01110000000","11111100010","00001100011","10000000001","01001010010","11000110000","00101111011","10100011001","01101001010","11100101000","00011101111","10010001101","01011011110","11010111100","00111110111","10110010101","01111000110","11110100100","00000010111","10001110101","01000100110","11001000100","00100001111","10101101101","01100111110","11101011100","00010011011","10011111001","01010101010","11011001000","00110000011","10111100001","01110110010","11111010000","00001010001","10000110011","01001100000","11000000010","00101001001","10100101011","01101111000","11100011010","00011011101","10010111111","01011101100","11010001110","00111000101","10110100111","01111110100","11110010110","00000110100","10001010110","01000000101","11001100111","00100101100","10101001110","01100011101","11101111111","00010111000","10011011010","01010001001","11011101011","00110100000","10111000010","01110010001","11111110011","00001110010","10000010000","01001000011","11000100001","00101101010","10100001000","01101011011","11100111001","00011111110","10010011100","01011001111","11010101101","00111100110","10110000100","01111010111","11110110101","00000001110","10001101100","01000111111","11001011101","00100010110","10101110100","01100100111","11101000101","00010000010","10011100000","01010110011","11011010001","00110011010","10111111000","01110101011","11111001001","00001001000","10000101010","01001111001","11000011011","00101010000","10100110010","01101100001","11100000011","00011000100","10010100110","01011110101","11010010111","00111011100","10110111110","01111101101","11110001111","00000101101","10001001111","01000011100","11001111110","00100110101","10101010111","01100000100","11101100110","00010100001","10011000011","01010010000","11011110010","00110111001","10111011011","01110001000","11111101010","00001101011","10000001001","01001011010","11000111000","00101110011","10100010001","01101000010","11100100000","00011100111","10010000101","01011010110","11010110100","00111111111","10110011101","01111001110","11110101100","00000011111","10001111101","01000101110","11001001100","00100000111","10101100101","01100110110","11101010100","00010010011","10011110001","01010100010","11011000000","00110001011","10111101001","01110111010","11111011000","00001011001","10000111011","01001101000","11000001010","00101000001","10100100011","01101110000","11100010010","00011010101","10010110111","01011100100","11010000110","00111001101","10110101111","01111111100","11110011110","00000111100","10001011110","01000001101","11001101111","00100100100","10101000110","01100010101","11101110111","00010110000","10011010010","01010000001","11011100011","00110101000","10111001010","01110011001","11111111011","00001111010","10000011000","01001001011","11000101001","00101100010","10100000000","01101010011","11100110001","00011110110","10010010100","01011000111","11010100101","00111101110","10110001100","01111011111","11110111101","00000000001","10001100011","01000110000","11001010010","00100011001","10101111011","01100101000","11101001010","00010001101","10011101111","01010111100","11011011110","00110010101","10111110111","01110100100","11111000110","00001000111","10000100101","01001110110","11000010100","00101011111","10100111101","01101101110","11100001100","00011001011","10010101001","01011111010","11010011000","00111010011","10110110001","01111100010","11110000000","00000100010","10001000000","01000010011","11001110001","00100111010","10101011000","01100001011","11101101001","00010101110","10011001100","01010011111","11011111101","00110110110","10111010100","01110000111","11111100101","00001100100","10000000110","01001010101","11000110111","00101111100","10100011110","01101001101","11100101111","00011101000","10010001010","01011011001","11010111011","00111110000","10110010010","01111000001","11110100011","00000010000","10001110010","01000100001","11001000011","00100001000","10101101010","01100111001","11101011011","00010011100","10011111110","01010101101","11011001111","00110000100","10111100110","01110110101","11111010111","00001010110","10000110100","01001100111","11000000101","00101001110","10100101100","01101111111","11100011101","00011011010","10010111000","01011101011","11010001001","00111000010","10110100000","01111110011","11110010001","00000110011","10001010001","01000000010","11001100000","00100101011","10101001001","01100011010","11101111000","00010111111","10011011101","01010001110","11011101100","00110100111","10111000101","01110010110","11111110100","00001110101","10000010111","01001000100","11000100110","00101101101","10100001111","01101011100","11100111110","00011111001","10010011011","01011001000","11010101010","00111100001","10110000011","01111010000","11110110010","00000001001","10001101011","01000111000","11001011010","00100010001","10101110011","01100100000","11101000010","00010000101","10011100111","01010110100","11011010110","00110011101","10111111111","01110101100","11111001110","00001001111","10000101101","01001111110","11000011100","00101010111","10100110101","01101100110","11100000100","00011000011","10010100001","01011110010","11010010000","00111011011","10110111001","01111101010","11110001000","00000101010","10001001000","01000011011","11001111001","00100110010","10101010000","01100000011","11101100001","00010100110","10011000100","01010010111","11011110101","00110111110","10111011100","01110001111","11111101101","00001101100","10000001110","01001011101","11000111111","00101110100","10100010110","01101000101","11100100111","00011100000","10010000010","01011010001","11010110011","00111111000","10110011010","01111001001","11110101011","00000011000","10001111010","01000101001","11001001011","00100000000","10101100010","01100110001","11101010011","00010010100","10011110110","01010100101","11011000111","00110001100","10111101110","01110111101","11111011111","00001011110","10000111100","01001101111","11000001101","00101000110","10100100100","01101110111","11100010101","00011010010","10010110000","01011100011","11010000001","00111001010","10110101000","01111111011","11110011001","00000111011","10001011001","01000001010","11001101000","00100100011","10101000001","01100010010","11101110000","00010110111","10011010101","01010000110","11011100100","00110101111","10111001101","01110011110","11111111100","00001111101","10000011111","01001001100","11000101110","00101100101","10100000111","01101010100","11100110110","00011110001","10010010011","01011000000","11010100010","00111101001","10110001011","01111011000","11110111010","00000000101","10001100111","01000110100","11001010110","00100011101","10101111111","01100101100","11101001110","00010001001","10011101011","01010111000","11011011010","00110010001","10111110011","01110100000","11111000010","00001000011","10000100001","01001110010","11000010000","00101011011","10100111001","01101101010","11100001000","00011001111","10010101101","01011111110","11010011100","00111010111","10110110101","01111100110","11110000100","00000100110","10001000100","01000010111","11001110101","00100111110","10101011100","01100001111","11101101101","00010101010","10011001000","01010011011","11011111001","00110110010","10111010000","01110000011","11111100001","00001100000","10000000010","01001010001","11000110011","00101111000","10100011010","01101001001","11100101011","00011101100","10010001110","01011011101","11010111111","00111110100","10110010110","01111000101","11110100111","00000010100","10001110110","01000100101","11001000111","00100001100","10101101110","01100111101","11101011111","00010011000","10011111010","01010101001","11011001011","00110000000","10111100010","01110110001","11111010011","00001010010","10000110000","01001100011","11000000001","00101001010","10100101000","01101111011","11100011001","00011011110","10010111100","01011101111","11010001101","00111000110","10110100100","01111110111","11110010101","00000110111","10001010101","01000000110","11001100100","00100101111","10101001101","01100011110","11101111100","00010111011","10011011001","01010001010","11011101000","00110100011","10111000001","01110010010","11111110000","00001110001","10000010011","01001000000","11000100010","00101101001","10100001011","01101011000","11100111010","00011111101","10010011111","01011001100","11010101110","00111100101","10110000111","01111010100","11110110110","00000001101","10001101111","01000111100","11001011110","00100010101","10101110111","01100100100","11101000110","00010000001","10011100011","01010110000","11011010010","00110011001","10111111011","01110101000","11111001010",
        "00001001011","10000101001","01001111010","11000011000","00101010011","10100110001","01101100010","11100000000","00011000111","10010100101","01011110110","11010010100","00111011111","10110111101","01111101110","11110001100","00000101110","10001001100","01000011111","11001111101","00100110110","10101010100","01100000111","11101100101","00010100010","10011000000","01010010011","11011110001","00110111010","10111011000","01110001011","11111101001","00001101000","10000001010","01001011001","11000111011","00101110000","10100010010","01101000001","11100100011","00011100100","10010000110","01011010101","11010110111","00111111100","10110011110","01111001101","11110101111","00000011100","10001111110","01000101101","11001001111","00100000100","10101100110","01100110101","11101010111","00010010000","10011110010","01010100001","11011000011","00110001000","10111101010","01110111001","11111011011","00001011010","10000111000","01001101011","11000001001","00101000010","10100100000","01101110011","11100010001","00011010110","10010110100","01011100111","11010000101","00111001110","10110101100","01111111111","11110011101","00000111111","10001011101","01000001110","11001101100","00100100111","10101000101","01100010110","11101110100","00010110011","10011010001","01010000010","11011100000","00110101011","10111001001","01110011010","11111111000","00001111001","10000011011","01001001000","11000101010","00101100001","10100000011","01101010000","11100110010","00011110101","10010010111","01011000100","11010100110","00111101101","10110001111","01111011100","11110111110","00000000011","10001100001","01000110010","11001010000","00100011011","10101111001","01100101010","11101001000","00010001111","10011101101","01010111110","11011011100","00110010111","10111110101","01110100110","11111000100","00001000101","10000100111","01001110100","11000010110","00101011101","10100111111","01101101100","11100001110","00011001001","10010101011","01011111000","11010011010","00111010001","10110110011","01111100000","11110000010","00000100000","10001000010","01000010001","11001110011","00100111000","10101011010","01100001001","11101101011","00010101100","10011001110","01010011101","11011111111","00110110100","10111010110","01110000101","11111100111","00001100110","10000000100","01001010111","11000110101","00101111110","10100011100","01101001111","11100101101","00011101010","10010001000","01011011011","11010111001","00111110010","10110010000","01111000011","11110100001","00000010010","10001110000","01000100011","11001000001","00100001010","10101101000","01100111011","11101011001","00010011110","10011111100","01010101111","11011001101","00110000110","10111100100","01110110111","11111010101","00001010100","10000110110","01001100101","11000000111","00101001100","10100101110","01101111101","11100011111","00011011000","10010111010","01011101001","11010001011","00111000000","10110100010","01111110001","11110010011","00000110001","10001010011","01000000000","11001100010","00100101001","10101001011","01100011000","11101111010","00010111101","10011011111","01010001100","11011101110","00110100101","10111000111","01110010100","11111110110","00001110111","10000010101","01001000110","11000100100","00101101111","10100001101","01101011110","11100111100","00011111011","10010011001","01011001010","11010101000","00111100011","10110000001","01111010010","11110110000","00000001011","10001101001","01000111010","11001011000","00100010011","10101110001","01100100010","11101000000","00010000111","10011100101","01010110110","11011010100","00110011111","10111111101","01110101110","11111001100","00001001101","10000101111","01001111100","11000011110","00101010101","10100110111","01101100100","11100000110","00011000001","10010100011","01011110000","11010010010","00111011001","10110111011","01111101000","11110001010","00000101000","10001001010","01000011001","11001111011","00100110000","10101010010","01100000001","11101100011","00010100100","10011000110","01010010101","11011110111","00110111100","10111011110","01110001101","11111101111","00001101110","10000001100","01001011111","11000111101","00101110110","10100010100","01101000111","11100100101","00011100010","10010000000","01011010011","11010110001","00111111010","10110011000","01111001011","11110101001","00000011010","10001111000","01000101011","11001001001","00100000010","10101100000","01100110011","11101010001","00010010110","10011110100","01010100111","11011000101","00110001110","10111101100","01110111111","11111011101","00001011100","10000111110","01001101101","11000001111","00101000100","10100100110","01101110101","11100010111","00011010000","10010110010","01011100001","11010000011","00111001000","10110101010","01111111001","11110011011","00000111001","10001011011","01000001000","11001101010","00100100001","10101000011","01100010000","11101110010","00010110101","10011010111","01010000100","11011100110","00110101101","10111001111","01110011100","11111111110","00001111111","10000011101","01001001110","11000101100","00101100111","10100000101","01101010110","11100110100","00011110011","10010010001","01011000010","11010100000","00111101011","10110001001","01111011010","11110111000","00000000111","10001100101","01000110110","11001010100","00100011111","10101111101","01100101110","11101001100","00010001011","10011101001","01010111010","11011011000","00110010011","10111110001","01110100010","11111000000","00001000001","10000100011","01001110000","11000010010","00101011001","10100111011","01101101000","11100001010","00011001101","10010101111","01011111100","11010011110","00111010101","10110110111","01111100100","11110000110","00000100100","10001000110","01000010101","11001110111","00100111100","10101011110","01100001101","11101101111","00010101000","10011001010","01010011001","11011111011","00110110000","10111010010","01110000001","11111100011","00001100010","10000000000","01001010011","11000110001","00101111010","10100011000","01101001011","11100101001","00011101110","10010001100","01011011111","11010111101","00111110110","10110010100","01111000111","11110100101","00000010110","10001110100","01000100111","11001000101","00100001110","10101101100","01100111111","11101011101","00010011010","10011111000","01010101011","11011001001","00110000010","10111100000","01110110011","11111010001","00001010000","10000110010","01001100001","11000000011","00101001000","10100101010","01101111001","11100011011","00011011100","10010111110","01011101101","11010001111","00111000100","10110100110","01111110101","11110010111","00000110101","10001010111","01000000100","11001100110","00100101101","10101001111","01100011100","11101111110","00010111001","10011011011","01010001000","11011101010","00110100001","10111000011","01110010000","11111110010","00001110011","10000010001","01001000010","11000100000","00101101011","10100001001","01101011010","11100111000","00011111111","10010011101","01011001110","11010101100","00111100111","10110000101","01111010110","11110110100","00000001111","10001101101","01000111110","11001011100","00100010111","10101110101","01100100110","11101000100","00010000011","10011100001","01010110010","11011010000","00110011011","10111111001","01110101010","11111001000","00001001001","10000101011","01001111000","11000011010","00101010001","10100110011","01101100000","11100000010","00011000101","10010100111","01011110100","11010010110","00111011101","10110111111","01111101100","11110001110","00000101100","10001001110","01000011101","11001111111","00100110100","10101010110","01100000101","11101100111","00010100000","10011000010","01010010001","11011110011","00110111000","10111011010","01110001001","11111101011","00001101010","10000001000","01001011011","11000111001","00101110010","10100010000","01101000011","11100100001","00011100110","10010000100","01011010111","11010110101","00111111110","10110011100","01111001111","11110101101","00000011110","10001111100","01000101111","11001001101","00100000110","10101100100","01100110111","11101010101","00010010010","10011110000","01010100011","11011000001","00110001010","10111101000","01110111011","11111011001","00001011000","10000111010","01001101001","11000001011","00101000000","10100100010","01101110001","11100010011","00011010100","10010110110","01011100101","11010000111","00111001100","10110101110","01111111101","11110011111","00000111101","10001011111","01000001100","11001101110","00100100101","10101000111","01100010100","11101110110","00010110001","10011010011","01010000000","11011100010","00110101001","10111001011","01110011000","11111111010","00001111011","10000011001","01001001010","11000101000","00101100011","10100000001","01101010010","11100110000","00011110111","10010010101","01011000110","11010100100","00111101111","10110001101","01111011110","11110111100");
        
      begin

      clk_tb <= (not(clk_tb) and end_sim) after T_CLK / 2;
      diff <= '1' when ((count="00000000000") and (output_expected /= outp)) else '0';
      
      output_expected <= outp_expected(t_integer);
      a_in_tb <= innp(0);

        test_CCG: CCG
        port map(
            clk => clk_tb,
            rst => rst_tb,
            a_in => a_in_tb,
            a_out => a_out_tb,
            c => c_out_tb
        );

        d_process: process(clk_tb, rst_tb) 
              begin
                if(rst_tb = '1') then
                  rst_tb <= '0' after T_RESET;
                elsif(rising_edge(clk_tb)) then
                      if(t_integer = 2047 and outp <= "00000000000")then end_sim <= '0';  end if;
                      if(count="000000000000") then
                          rst_tb <= '1'; 
                          t_integer <= (t_integer + 1); 
                          count <= "110000000000";
                          innp <= std_logic_vector(to_unsigned(t_integer+1, innp'length));
                          outp <= "00000000000";
                      else
                          count <= '0' & count(11 downto 1) ;
                          innp <= '0' & innp(10 downto 1) ;
                          outp <= outp(9 downto 0) & c_out_tb ;                          
                      end if;
                end if;
              end process;
    end bench;
